`timescale 1ns / 1ps
module Sliding_average_filter#(
    parameter WINDOW_WIDTH = 10,//窗口位宽
    parameter en_sample_interval = 0,//使能采样间隔
    parameter DATA_WIDTH = 16  //数据位宽
)(
    input clk,
    input [DATA_WIDTH-1:0]i_data,
    input i_valid,
    input [7:0]i_sample_interval,
    output [DATA_WIDTH-1:0]o_data,
    output o_valid
    );
localparam WINDOW_LENGTH = 2**WINDOW_WIDTH;
//--------------------------------------------------------
//   256级寄存器移位缓存数据
//--------------------------------------------------------
reg [DATA_WIDTH-1:0] din_reg [WINDOW_LENGTH-1:0];
integer j; 
//采样
reg [7:0]samp_cnt=0;
reg [DATA_WIDTH-1:0]r_data;
reg r_valid;
always @(posedge clk) begin
    if(en_sample_interval)begin
        if(i_valid)begin
            if(samp_cnt>=i_sample_interval-1)begin
                samp_cnt<=0;
                r_data<=i_data;
            end
            else begin
                samp_cnt<=samp_cnt+1;
            end
        end
        r_valid<=(i_valid & samp_cnt==i_sample_interval-1) ? 1:0;
    end
    else begin
        if(i_valid)begin
            r_data<=i_data;
            r_valid<=1;
        end
        else r_valid<=0;
    end
end
always @ (posedge clk)
begin
    if(r_valid)begin
        din_reg[0] <= r_data;
        for (j=0; j<WINDOW_LENGTH-1; j=j+1)
            din_reg[j+1] <= din_reg[j];
    end
end

//--------------------------------------------------------
//   计算基带信号连续256个数据的均值
//--------------------------------------------------------    
reg signed [DATA_WIDTH+WINDOW_WIDTH-1:0] sum;
always @ (posedge clk)begin
    if(r_valid)begin
        //将最老的数据换为最新的数据
        sum <= sum + {{(WINDOW_WIDTH){r_data[DATA_WIDTH-1]}},r_data} 
                    - {{(WINDOW_WIDTH){din_reg[WINDOW_LENGTH-1][DATA_WIDTH-1]}},din_reg[WINDOW_LENGTH-1]};   
    end
end
assign o_data = sum[DATA_WIDTH+WINDOW_WIDTH-1:WINDOW_WIDTH];  //右移8bit等效为÷256    
assign o_valid = r_valid;
endmodule
